library verilog;
use verilog.vl_types.all;
entity bcd_coder_vlg_check_tst is
    port(
        yout            : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end bcd_coder_vlg_check_tst;
