library verilog;
use verilog.vl_types.all;
entity bin2bcd_vlg_vec_tst is
end bin2bcd_vlg_vec_tst;
